\+---doing_so_inst1: doing_so
    --- CLK_FREQ    => 10,
    --- SCL_FREQ    => 4
    --- Reset_s          =>   Reset_s,
    --- Clk_4MHz         =>   Clk_4MHz,
    --- Signal_in        =>   sig_internal,
    --- Signal_out       =>   sig_out,
    --- Signal_open      =>   open

\+---doing_so_inst2: doing_so
    --- Reset_s      =>Reset_s,
    --- Clk_4MHz     =>Clk_100MHz,
    --- Signal_in    =>sig_internal,
    --- Signal_out   =>open,
    --- Signal_open  =>open

\+---doing_so_inst3: doing_so
    --- 72
    --- 10
    --- Reset_s
    --- Clk_120MHz
    --- sig_internal
    --- sig_out2
    --- open

\+---doing_so_inst4: doing_so
    --- Reset_s      =>Reset_s,
    --- Clk_4MHz     =>Clk_100MHz,
    --- Signal_in    =>sig_internal,
    --- Signal_out   =>open,
    --- Signal_open  =>open